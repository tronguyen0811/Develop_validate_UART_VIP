interface uart_if();

  logic tx;
  logic rx;
  
endinterface
